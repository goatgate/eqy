// This is the unpowered netlist.
module spm (clk,
p,
rst,
y,
x);
input clk;
output p;
input rst;
input y;
input [31:0] x;

wire _000_;
wire _001_;
wire _002_;
wire _003_;
wire _004_;
wire _005_;
wire _006_;
wire _007_;
wire _008_;
wire _009_;
wire _010_;
wire _011_;
wire _012_;
wire _013_;
wire _014_;
wire _015_;
wire _016_;
wire _017_;
wire _018_;
wire _019_;
wire _020_;
wire _021_;
wire _022_;
wire _023_;
wire _024_;
wire _025_;
wire _026_;
wire _027_;
wire _028_;
wire _029_;
wire _030_;
wire _031_;
wire _032_;
wire _033_;
wire _034_;
wire _035_;
wire _036_;
wire _037_;
wire _038_;
wire _039_;
wire _040_;
wire _041_;
wire _042_;
wire _043_;
wire _044_;
wire _045_;
wire _046_;
wire _047_;
wire _048_;
wire _049_;
wire _050_;
wire _051_;
wire _052_;
wire _053_;
wire _054_;
wire _055_;
wire _056_;
wire _057_;
wire _058_;
wire _059_;
wire _060_;
wire _061_;
wire _062_;
wire _063_;
wire _064_;
wire _065_;
wire _066_;
wire _067_;
wire _068_;
wire _069_;
wire _070_;
wire _071_;
wire _072_;
wire _073_;
wire _074_;
wire _075_;
wire _076_;
wire _077_;
wire _078_;
wire _079_;
wire _080_;
wire _081_;
wire _082_;
wire _083_;
wire _084_;
wire _085_;
wire _086_;
wire _087_;
wire _088_;
wire _089_;
wire _090_;
wire _091_;
wire _092_;
wire _093_;
wire _094_;
wire _095_;
wire _096_;
wire _097_;
wire _098_;
wire _099_;
wire _100_;
wire _101_;
wire _102_;
wire _103_;
wire _104_;
wire _105_;
wire _106_;
wire _107_;
wire _108_;
wire _109_;
wire _110_;
wire _111_;
wire _112_;
wire _113_;
wire _114_;
wire _115_;
wire _116_;
wire _117_;
wire _118_;
wire _119_;
wire _120_;
wire _121_;
wire _122_;
wire _123_;
wire _124_;
wire _125_;
wire _126_;
wire _127_;
wire _128_;
wire _129_;
wire _130_;
wire _131_;
wire _132_;
wire _133_;
wire _134_;
wire _135_;
wire _136_;
wire _137_;
wire _138_;
wire _139_;
wire _140_;
wire _141_;
wire _142_;
wire _143_;
wire _144_;
wire _145_;
wire _146_;
wire _147_;
wire _148_;
wire _149_;
wire _150_;
wire _151_;
wire _152_;
wire _153_;
wire _154_;
wire _155_;
wire _156_;
wire _157_;
wire _158_;
wire _159_;
wire _160_;
wire _161_;
wire _162_;
wire _163_;
wire _164_;
wire _165_;
wire _166_;
wire _167_;
wire _168_;
wire _169_;
wire _170_;
wire _171_;
wire _172_;
wire _173_;
wire _174_;
wire _175_;
wire _176_;
wire _177_;
wire _178_;
wire _179_;
wire _180_;
wire _181_;
wire _182_;
wire _183_;
wire _184_;
wire _185_;
wire _186_;
wire _187_;
wire _188_;
wire _189_;
wire _190_;
wire _191_;
wire _192_;
wire _193_;
wire _194_;
wire _195_;
wire _196_;
wire _197_;
wire _198_;
wire _199_;
wire _200_;
wire _201_;
wire _202_;
wire _203_;
wire _204_;
wire _205_;
wire clknet_0_clk;
wire clknet_3_0__leaf_clk;
wire clknet_3_1__leaf_clk;
wire clknet_3_2__leaf_clk;
wire clknet_3_3__leaf_clk;
wire clknet_3_4__leaf_clk;
wire clknet_3_5__leaf_clk;
wire clknet_3_6__leaf_clk;
wire clknet_3_7__leaf_clk;
wire \csa0.hsum2 ;
wire \csa0.sc ;
wire \csa0.y ;
wire \genblk1[10].csa.hsum2 ;
wire \genblk1[10].csa.sc ;
wire \genblk1[10].csa.sum ;
wire \genblk1[10].csa.y ;
wire \genblk1[11].csa.hsum2 ;
wire \genblk1[11].csa.sc ;
wire \genblk1[11].csa.y ;
wire \genblk1[12].csa.hsum2 ;
wire \genblk1[12].csa.sc ;
wire \genblk1[12].csa.y ;
wire \genblk1[13].csa.hsum2 ;
wire \genblk1[13].csa.sc ;
wire \genblk1[13].csa.y ;
wire \genblk1[14].csa.hsum2 ;
wire \genblk1[14].csa.sc ;
wire \genblk1[14].csa.y ;
wire \genblk1[15].csa.hsum2 ;
wire \genblk1[15].csa.sc ;
wire \genblk1[15].csa.y ;
wire \genblk1[16].csa.hsum2 ;
wire \genblk1[16].csa.sc ;
wire \genblk1[16].csa.y ;
wire \genblk1[17].csa.hsum2 ;
wire \genblk1[17].csa.sc ;
wire \genblk1[17].csa.y ;
wire \genblk1[18].csa.hsum2 ;
wire \genblk1[18].csa.sc ;
wire \genblk1[18].csa.y ;
wire \genblk1[19].csa.hsum2 ;
wire \genblk1[19].csa.sc ;
wire \genblk1[19].csa.y ;
wire \genblk1[1].csa.hsum2 ;
wire \genblk1[1].csa.sc ;
wire \genblk1[1].csa.y ;
wire \genblk1[20].csa.hsum2 ;
wire \genblk1[20].csa.sc ;
wire \genblk1[20].csa.y ;
wire \genblk1[21].csa.hsum2 ;
wire \genblk1[21].csa.sc ;
wire \genblk1[21].csa.y ;
wire \genblk1[22].csa.hsum2 ;
wire \genblk1[22].csa.sc ;
wire \genblk1[22].csa.y ;
wire \genblk1[23].csa.hsum2 ;
wire \genblk1[23].csa.sc ;
wire \genblk1[23].csa.y ;
wire \genblk1[24].csa.hsum2 ;
wire \genblk1[24].csa.sc ;
wire \genblk1[24].csa.y ;
wire \genblk1[25].csa.hsum2 ;
wire \genblk1[25].csa.sc ;
wire \genblk1[25].csa.y ;
wire \genblk1[26].csa.hsum2 ;
wire \genblk1[26].csa.sc ;
wire \genblk1[26].csa.y ;
wire \genblk1[27].csa.hsum2 ;
wire \genblk1[27].csa.sc ;
wire \genblk1[27].csa.y ;
wire \genblk1[28].csa.hsum2 ;
wire \genblk1[28].csa.sc ;
wire \genblk1[28].csa.y ;
wire \genblk1[29].csa.hsum2 ;
wire \genblk1[29].csa.sc ;
wire \genblk1[29].csa.y ;
wire \genblk1[2].csa.hsum2 ;
wire \genblk1[2].csa.sc ;
wire \genblk1[2].csa.y ;
wire \genblk1[30].csa.hsum2 ;
wire \genblk1[30].csa.sc ;
wire \genblk1[30].csa.y ;
wire \genblk1[3].csa.hsum2 ;
wire \genblk1[3].csa.sc ;
wire \genblk1[3].csa.y ;
wire \genblk1[4].csa.hsum2 ;
wire \genblk1[4].csa.sc ;
wire \genblk1[4].csa.y ;
wire \genblk1[5].csa.hsum2 ;
wire \genblk1[5].csa.sc ;
wire \genblk1[5].csa.y ;
wire \genblk1[6].csa.hsum2 ;
wire \genblk1[6].csa.sc ;
wire \genblk1[6].csa.y ;
wire \genblk1[7].csa.hsum2 ;
wire \genblk1[7].csa.sc ;
wire \genblk1[7].csa.y ;
wire \genblk1[8].csa.hsum2 ;
wire \genblk1[8].csa.sc ;
wire \genblk1[8].csa.y ;
wire \genblk1[9].csa.hsum2 ;
wire \genblk1[9].csa.sc ;
wire net1;
wire net10;
wire net11;
wire net12;
wire net13;
wire net14;
wire net15;
wire net16;
wire net17;
wire net18;
wire net19;
wire net2;
wire net20;
wire net21;
wire net22;
wire net23;
wire net24;
wire net25;
wire net26;
wire net27;
wire net28;
wire net29;
wire net3;
wire net30;
wire net31;
wire net32;
wire net33;
wire net34;
wire net35;
wire net4;
wire net5;
wire net6;
wire net7;
wire net8;
wire net9;
wire \tcmp.z ;

sky130_fd_sc_hd__decap_8 FILLER_0_102 ();
sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
sky130_fd_sc_hd__decap_12 FILLER_0_113 ();
sky130_fd_sc_hd__decap_6 FILLER_0_125 ();
sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
sky130_fd_sc_hd__decap_8 FILLER_0_141 ();
sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
sky130_fd_sc_hd__decap_12 FILLER_0_15 ();
sky130_fd_sc_hd__decap_4 FILLER_0_153 ();
sky130_fd_sc_hd__decap_4 FILLER_0_164 ();
sky130_fd_sc_hd__decap_4 FILLER_0_169 ();
sky130_fd_sc_hd__fill_1 FILLER_0_173 ();
sky130_fd_sc_hd__decap_6 FILLER_0_177 ();
sky130_fd_sc_hd__fill_1 FILLER_0_183 ();
sky130_fd_sc_hd__decap_6 FILLER_0_187 ();
sky130_fd_sc_hd__fill_1 FILLER_0_193 ();
sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
sky130_fd_sc_hd__decap_12 FILLER_0_29 ();
sky130_fd_sc_hd__decap_12 FILLER_0_3 ();
sky130_fd_sc_hd__decap_12 FILLER_0_41 ();
sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
sky130_fd_sc_hd__decap_12 FILLER_0_57 ();
sky130_fd_sc_hd__decap_12 FILLER_0_69 ();
sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
sky130_fd_sc_hd__decap_12 FILLER_0_85 ();
sky130_fd_sc_hd__fill_2 FILLER_0_97 ();
sky130_fd_sc_hd__decap_4 FILLER_10_113 ();
sky130_fd_sc_hd__decap_3 FILLER_10_137 ();
sky130_fd_sc_hd__decap_8 FILLER_10_141 ();
sky130_fd_sc_hd__fill_2 FILLER_10_149 ();
sky130_fd_sc_hd__decap_12 FILLER_10_15 ();
sky130_fd_sc_hd__decap_8 FILLER_10_171 ();
sky130_fd_sc_hd__decap_4 FILLER_10_182 ();
sky130_fd_sc_hd__decap_4 FILLER_10_189 ();
sky130_fd_sc_hd__fill_1 FILLER_10_193 ();
sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
sky130_fd_sc_hd__decap_8 FILLER_10_29 ();
sky130_fd_sc_hd__decap_12 FILLER_10_3 ();
sky130_fd_sc_hd__fill_1 FILLER_10_37 ();
sky130_fd_sc_hd__decap_4 FILLER_10_58 ();
sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
sky130_fd_sc_hd__decap_8 FILLER_10_85 ();
sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
sky130_fd_sc_hd__decap_8 FILLER_11_113 ();
sky130_fd_sc_hd__decap_4 FILLER_11_12 ();
sky130_fd_sc_hd__fill_2 FILLER_11_121 ();
sky130_fd_sc_hd__decap_12 FILLER_11_143 ();
sky130_fd_sc_hd__decap_12 FILLER_11_155 ();
sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
sky130_fd_sc_hd__decap_3 FILLER_11_191 ();
sky130_fd_sc_hd__decap_4 FILLER_11_21 ();
sky130_fd_sc_hd__decap_6 FILLER_11_28 ();
sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
sky130_fd_sc_hd__decap_4 FILLER_11_57 ();
sky130_fd_sc_hd__decap_8 FILLER_11_81 ();
sky130_fd_sc_hd__fill_1 FILLER_11_89 ();
sky130_fd_sc_hd__fill_1 FILLER_12_105 ();
sky130_fd_sc_hd__decap_12 FILLER_12_126 ();
sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
sky130_fd_sc_hd__decap_8 FILLER_12_163 ();
sky130_fd_sc_hd__decap_3 FILLER_12_191 ();
sky130_fd_sc_hd__decap_6 FILLER_12_22 ();
sky130_fd_sc_hd__decap_4 FILLER_12_29 ();
sky130_fd_sc_hd__decap_12 FILLER_12_3 ();
sky130_fd_sc_hd__decap_8 FILLER_12_53 ();
sky130_fd_sc_hd__fill_1 FILLER_12_61 ();
sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
sky130_fd_sc_hd__decap_12 FILLER_12_85 ();
sky130_fd_sc_hd__decap_8 FILLER_12_97 ();
sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
sky130_fd_sc_hd__decap_12 FILLER_13_113 ();
sky130_fd_sc_hd__decap_12 FILLER_13_125 ();
sky130_fd_sc_hd__decap_12 FILLER_13_137 ();
sky130_fd_sc_hd__decap_12 FILLER_13_149 ();
sky130_fd_sc_hd__decap_4 FILLER_13_16 ();
sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
sky130_fd_sc_hd__decap_3 FILLER_13_169 ();
sky130_fd_sc_hd__fill_2 FILLER_13_192 ();
sky130_fd_sc_hd__fill_1 FILLER_13_20 ();
sky130_fd_sc_hd__decap_8 FILLER_13_24 ();
sky130_fd_sc_hd__decap_6 FILLER_13_3 ();
sky130_fd_sc_hd__fill_2 FILLER_13_32 ();
sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
sky130_fd_sc_hd__decap_12 FILLER_13_57 ();
sky130_fd_sc_hd__decap_4 FILLER_13_69 ();
sky130_fd_sc_hd__decap_12 FILLER_13_93 ();
sky130_fd_sc_hd__fill_1 FILLER_14_11 ();
sky130_fd_sc_hd__decap_4 FILLER_14_113 ();
sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
sky130_fd_sc_hd__decap_4 FILLER_14_15 ();
sky130_fd_sc_hd__decap_4 FILLER_14_163 ();
sky130_fd_sc_hd__decap_6 FILLER_14_187 ();
sky130_fd_sc_hd__fill_1 FILLER_14_193 ();
sky130_fd_sc_hd__decap_6 FILLER_14_22 ();
sky130_fd_sc_hd__decap_4 FILLER_14_29 ();
sky130_fd_sc_hd__decap_8 FILLER_14_3 ();
sky130_fd_sc_hd__decap_4 FILLER_14_53 ();
sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
sky130_fd_sc_hd__decap_8 FILLER_14_85 ();
sky130_fd_sc_hd__decap_4 FILLER_15_108 ();
sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
sky130_fd_sc_hd__decap_4 FILLER_15_135 ();
sky130_fd_sc_hd__decap_8 FILLER_15_159 ();
sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
sky130_fd_sc_hd__decap_4 FILLER_15_18 ();
sky130_fd_sc_hd__decap_3 FILLER_15_191 ();
sky130_fd_sc_hd__decap_8 FILLER_15_25 ();
sky130_fd_sc_hd__decap_3 FILLER_15_3 ();
sky130_fd_sc_hd__fill_1 FILLER_15_33 ();
sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
sky130_fd_sc_hd__decap_12 FILLER_15_57 ();
sky130_fd_sc_hd__decap_6 FILLER_15_69 ();
sky130_fd_sc_hd__fill_1 FILLER_15_75 ();
sky130_fd_sc_hd__decap_4 FILLER_15_9 ();
sky130_fd_sc_hd__decap_12 FILLER_15_96 ();
sky130_fd_sc_hd__decap_12 FILLER_16_109 ();
sky130_fd_sc_hd__decap_3 FILLER_16_11 ();
sky130_fd_sc_hd__decap_12 FILLER_16_121 ();
sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
sky130_fd_sc_hd__decap_4 FILLER_16_163 ();
sky130_fd_sc_hd__decap_6 FILLER_16_187 ();
sky130_fd_sc_hd__fill_1 FILLER_16_193 ();
sky130_fd_sc_hd__decap_6 FILLER_16_21 ();
sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
sky130_fd_sc_hd__decap_4 FILLER_16_29 ();
sky130_fd_sc_hd__decap_8 FILLER_16_3 ();
sky130_fd_sc_hd__decap_8 FILLER_16_53 ();
sky130_fd_sc_hd__fill_1 FILLER_16_61 ();
sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
sky130_fd_sc_hd__decap_12 FILLER_16_85 ();
sky130_fd_sc_hd__decap_12 FILLER_16_97 ();
sky130_fd_sc_hd__decap_6 FILLER_17_106 ();
sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
sky130_fd_sc_hd__decap_8 FILLER_17_12 ();
sky130_fd_sc_hd__decap_12 FILLER_17_135 ();
sky130_fd_sc_hd__decap_12 FILLER_17_147 ();
sky130_fd_sc_hd__decap_8 FILLER_17_159 ();
sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
sky130_fd_sc_hd__decap_12 FILLER_17_174 ();
sky130_fd_sc_hd__decap_8 FILLER_17_186 ();
sky130_fd_sc_hd__fill_1 FILLER_17_20 ();
sky130_fd_sc_hd__decap_8 FILLER_17_24 ();
sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
sky130_fd_sc_hd__fill_1 FILLER_17_32 ();
sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
sky130_fd_sc_hd__decap_12 FILLER_17_57 ();
sky130_fd_sc_hd__decap_12 FILLER_17_69 ();
sky130_fd_sc_hd__decap_4 FILLER_17_81 ();
sky130_fd_sc_hd__fill_1 FILLER_17_85 ();
sky130_fd_sc_hd__decap_12 FILLER_18_116 ();
sky130_fd_sc_hd__decap_12 FILLER_18_128 ();
sky130_fd_sc_hd__decap_12 FILLER_18_14 ();
sky130_fd_sc_hd__decap_12 FILLER_18_141 ();
sky130_fd_sc_hd__decap_4 FILLER_18_153 ();
sky130_fd_sc_hd__decap_12 FILLER_18_177 ();
sky130_fd_sc_hd__decap_4 FILLER_18_189 ();
sky130_fd_sc_hd__fill_1 FILLER_18_193 ();
sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
sky130_fd_sc_hd__decap_4 FILLER_18_29 ();
sky130_fd_sc_hd__decap_4 FILLER_18_3 ();
sky130_fd_sc_hd__decap_12 FILLER_18_53 ();
sky130_fd_sc_hd__decap_12 FILLER_18_65 ();
sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
sky130_fd_sc_hd__decap_8 FILLER_18_85 ();
sky130_fd_sc_hd__decap_3 FILLER_18_93 ();
sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
sky130_fd_sc_hd__decap_6 FILLER_19_113 ();
sky130_fd_sc_hd__decap_4 FILLER_19_12 ();
sky130_fd_sc_hd__decap_4 FILLER_19_139 ();
sky130_fd_sc_hd__decap_4 FILLER_19_163 ();
sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
sky130_fd_sc_hd__decap_3 FILLER_19_169 ();
sky130_fd_sc_hd__decap_12 FILLER_19_19 ();
sky130_fd_sc_hd__fill_2 FILLER_19_192 ();
sky130_fd_sc_hd__decap_6 FILLER_19_3 ();
sky130_fd_sc_hd__fill_2 FILLER_19_31 ();
sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
sky130_fd_sc_hd__decap_6 FILLER_19_57 ();
sky130_fd_sc_hd__decap_6 FILLER_19_83 ();
sky130_fd_sc_hd__fill_1 FILLER_19_89 ();
sky130_fd_sc_hd__decap_3 FILLER_1_109 ();
sky130_fd_sc_hd__decap_3 FILLER_1_113 ();
sky130_fd_sc_hd__decap_12 FILLER_1_119 ();
sky130_fd_sc_hd__fill_1 FILLER_1_131 ();
sky130_fd_sc_hd__decap_12 FILLER_1_139 ();
sky130_fd_sc_hd__decap_12 FILLER_1_15 ();
sky130_fd_sc_hd__decap_4 FILLER_1_158 ();
sky130_fd_sc_hd__fill_1 FILLER_1_162 ();
sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
sky130_fd_sc_hd__decap_4 FILLER_1_169 ();
sky130_fd_sc_hd__fill_1 FILLER_1_173 ();
sky130_fd_sc_hd__decap_4 FILLER_1_181 ();
sky130_fd_sc_hd__decap_4 FILLER_1_190 ();
sky130_fd_sc_hd__decap_12 FILLER_1_27 ();
sky130_fd_sc_hd__decap_12 FILLER_1_3 ();
sky130_fd_sc_hd__decap_6 FILLER_1_39 ();
sky130_fd_sc_hd__fill_1 FILLER_1_45 ();
sky130_fd_sc_hd__decap_6 FILLER_1_49 ();
sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
sky130_fd_sc_hd__decap_6 FILLER_1_57 ();
sky130_fd_sc_hd__fill_1 FILLER_1_63 ();
sky130_fd_sc_hd__decap_8 FILLER_1_71 ();
sky130_fd_sc_hd__fill_1 FILLER_1_79 ();
sky130_fd_sc_hd__decap_4 FILLER_1_87 ();
sky130_fd_sc_hd__decap_12 FILLER_1_97 ();
sky130_fd_sc_hd__decap_8 FILLER_20_129 ();
sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
sky130_fd_sc_hd__fill_1 FILLER_20_15 ();
sky130_fd_sc_hd__decap_4 FILLER_20_163 ();
sky130_fd_sc_hd__decap_6 FILLER_20_187 ();
sky130_fd_sc_hd__fill_1 FILLER_20_193 ();
sky130_fd_sc_hd__decap_6 FILLER_20_22 ();
sky130_fd_sc_hd__decap_4 FILLER_20_29 ();
sky130_fd_sc_hd__decap_12 FILLER_20_3 ();
sky130_fd_sc_hd__decap_8 FILLER_20_53 ();
sky130_fd_sc_hd__fill_1 FILLER_20_61 ();
sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
sky130_fd_sc_hd__decap_12 FILLER_20_85 ();
sky130_fd_sc_hd__decap_12 FILLER_20_97 ();
sky130_fd_sc_hd__decap_8 FILLER_21_103 ();
sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
sky130_fd_sc_hd__decap_6 FILLER_21_113 ();
sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
sky130_fd_sc_hd__decap_4 FILLER_21_12 ();
sky130_fd_sc_hd__decap_12 FILLER_21_140 ();
sky130_fd_sc_hd__decap_12 FILLER_21_152 ();
sky130_fd_sc_hd__decap_4 FILLER_21_164 ();
sky130_fd_sc_hd__decap_3 FILLER_21_169 ();
sky130_fd_sc_hd__fill_2 FILLER_21_192 ();
sky130_fd_sc_hd__decap_4 FILLER_21_21 ();
sky130_fd_sc_hd__decap_4 FILLER_21_28 ();
sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
sky130_fd_sc_hd__fill_1 FILLER_21_32 ();
sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
sky130_fd_sc_hd__decap_4 FILLER_21_79 ();
sky130_fd_sc_hd__decap_12 FILLER_22_109 ();
sky130_fd_sc_hd__decap_12 FILLER_22_121 ();
sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
sky130_fd_sc_hd__decap_12 FILLER_22_146 ();
sky130_fd_sc_hd__fill_1 FILLER_22_15 ();
sky130_fd_sc_hd__decap_12 FILLER_22_158 ();
sky130_fd_sc_hd__decap_12 FILLER_22_170 ();
sky130_fd_sc_hd__decap_4 FILLER_22_182 ();
sky130_fd_sc_hd__decap_4 FILLER_22_189 ();
sky130_fd_sc_hd__decap_4 FILLER_22_19 ();
sky130_fd_sc_hd__fill_1 FILLER_22_193 ();
sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
sky130_fd_sc_hd__decap_12 FILLER_22_29 ();
sky130_fd_sc_hd__decap_12 FILLER_22_3 ();
sky130_fd_sc_hd__decap_12 FILLER_22_41 ();
sky130_fd_sc_hd__fill_1 FILLER_22_53 ();
sky130_fd_sc_hd__decap_8 FILLER_22_74 ();
sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
sky130_fd_sc_hd__decap_12 FILLER_22_85 ();
sky130_fd_sc_hd__decap_12 FILLER_22_97 ();
sky130_fd_sc_hd__decap_4 FILLER_23_103 ();
sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
sky130_fd_sc_hd__decap_8 FILLER_23_118 ();
sky130_fd_sc_hd__decap_12 FILLER_23_12 ();
sky130_fd_sc_hd__decap_4 FILLER_23_129 ();
sky130_fd_sc_hd__decap_4 FILLER_23_136 ();
sky130_fd_sc_hd__decap_4 FILLER_23_143 ();
sky130_fd_sc_hd__decap_4 FILLER_23_150 ();
sky130_fd_sc_hd__decap_4 FILLER_23_157 ();
sky130_fd_sc_hd__decap_4 FILLER_23_164 ();
sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
sky130_fd_sc_hd__decap_8 FILLER_23_174 ();
sky130_fd_sc_hd__fill_2 FILLER_23_182 ();
sky130_fd_sc_hd__decap_6 FILLER_23_187 ();
sky130_fd_sc_hd__fill_1 FILLER_23_193 ();
sky130_fd_sc_hd__decap_12 FILLER_23_24 ();
sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
sky130_fd_sc_hd__decap_12 FILLER_23_36 ();
sky130_fd_sc_hd__decap_8 FILLER_23_48 ();
sky130_fd_sc_hd__decap_12 FILLER_23_57 ();
sky130_fd_sc_hd__decap_3 FILLER_23_69 ();
sky130_fd_sc_hd__decap_12 FILLER_23_75 ();
sky130_fd_sc_hd__decap_6 FILLER_23_87 ();
sky130_fd_sc_hd__decap_4 FILLER_23_96 ();
sky130_fd_sc_hd__decap_4 FILLER_24_103 ();
sky130_fd_sc_hd__decap_4 FILLER_24_110 ();
sky130_fd_sc_hd__decap_4 FILLER_24_120 ();
sky130_fd_sc_hd__decap_6 FILLER_24_127 ();
sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
sky130_fd_sc_hd__decap_6 FILLER_24_149 ();
sky130_fd_sc_hd__decap_4 FILLER_24_162 ();
sky130_fd_sc_hd__decap_12 FILLER_24_169 ();
sky130_fd_sc_hd__fill_1 FILLER_24_181 ();
sky130_fd_sc_hd__decap_4 FILLER_24_189 ();
sky130_fd_sc_hd__fill_1 FILLER_24_193 ();
sky130_fd_sc_hd__decap_6 FILLER_24_22 ();
sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
sky130_fd_sc_hd__decap_3 FILLER_24_3 ();
sky130_fd_sc_hd__decap_6 FILLER_24_36 ();
sky130_fd_sc_hd__decap_8 FILLER_24_49 ();
sky130_fd_sc_hd__fill_2 FILLER_24_57 ();
sky130_fd_sc_hd__decap_4 FILLER_24_62 ();
sky130_fd_sc_hd__decap_4 FILLER_24_69 ();
sky130_fd_sc_hd__decap_6 FILLER_24_78 ();
sky130_fd_sc_hd__decap_4 FILLER_24_85 ();
sky130_fd_sc_hd__decap_6 FILLER_24_9 ();
sky130_fd_sc_hd__decap_4 FILLER_24_96 ();
sky130_fd_sc_hd__decap_4 FILLER_25_107 ();
sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
sky130_fd_sc_hd__decap_4 FILLER_25_122 ();
sky130_fd_sc_hd__decap_4 FILLER_25_133 ();
sky130_fd_sc_hd__decap_8 FILLER_25_143 ();
sky130_fd_sc_hd__fill_1 FILLER_25_151 ();
sky130_fd_sc_hd__decap_8 FILLER_25_159 ();
sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
sky130_fd_sc_hd__decap_4 FILLER_25_178 ();
sky130_fd_sc_hd__decap_4 FILLER_25_189 ();
sky130_fd_sc_hd__decap_4 FILLER_25_19 ();
sky130_fd_sc_hd__fill_1 FILLER_25_193 ();
sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
sky130_fd_sc_hd__decap_4 FILLER_25_30 ();
sky130_fd_sc_hd__decap_4 FILLER_25_41 ();
sky130_fd_sc_hd__decap_4 FILLER_25_52 ();
sky130_fd_sc_hd__decap_6 FILLER_25_57 ();
sky130_fd_sc_hd__decap_4 FILLER_25_70 ();
sky130_fd_sc_hd__decap_4 FILLER_25_8 ();
sky130_fd_sc_hd__decap_8 FILLER_25_81 ();
sky130_fd_sc_hd__fill_2 FILLER_25_89 ();
sky130_fd_sc_hd__decap_4 FILLER_25_98 ();
sky130_fd_sc_hd__decap_12 FILLER_26_105 ();
sky130_fd_sc_hd__decap_3 FILLER_26_117 ();
sky130_fd_sc_hd__decap_12 FILLER_26_125 ();
sky130_fd_sc_hd__decap_3 FILLER_26_137 ();
sky130_fd_sc_hd__decap_4 FILLER_26_14 ();
sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
sky130_fd_sc_hd__decap_8 FILLER_26_147 ();
sky130_fd_sc_hd__fill_2 FILLER_26_155 ();
sky130_fd_sc_hd__decap_6 FILLER_26_162 ();
sky130_fd_sc_hd__fill_1 FILLER_26_168 ();
sky130_fd_sc_hd__decap_4 FILLER_26_172 ();
sky130_fd_sc_hd__decap_6 FILLER_26_179 ();
sky130_fd_sc_hd__decap_4 FILLER_26_190 ();
sky130_fd_sc_hd__decap_6 FILLER_26_22 ();
sky130_fd_sc_hd__decap_12 FILLER_26_29 ();
sky130_fd_sc_hd__decap_4 FILLER_26_3 ();
sky130_fd_sc_hd__decap_8 FILLER_26_41 ();
sky130_fd_sc_hd__decap_8 FILLER_26_54 ();
sky130_fd_sc_hd__fill_2 FILLER_26_62 ();
sky130_fd_sc_hd__decap_4 FILLER_26_67 ();
sky130_fd_sc_hd__fill_1 FILLER_26_7 ();
sky130_fd_sc_hd__fill_1 FILLER_26_71 ();
sky130_fd_sc_hd__decap_4 FILLER_26_75 ();
sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
sky130_fd_sc_hd__decap_12 FILLER_26_93 ();
sky130_fd_sc_hd__decap_8 FILLER_27_101 ();
sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
sky130_fd_sc_hd__decap_12 FILLER_27_118 ();
sky130_fd_sc_hd__decap_4 FILLER_27_13 ();
sky130_fd_sc_hd__fill_1 FILLER_27_130 ();
sky130_fd_sc_hd__decap_4 FILLER_27_138 ();
sky130_fd_sc_hd__decap_8 FILLER_27_145 ();
sky130_fd_sc_hd__fill_2 FILLER_27_153 ();
sky130_fd_sc_hd__decap_4 FILLER_27_158 ();
sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
sky130_fd_sc_hd__decap_6 FILLER_27_174 ();
sky130_fd_sc_hd__decap_4 FILLER_27_185 ();
sky130_fd_sc_hd__fill_2 FILLER_27_192 ();
sky130_fd_sc_hd__decap_4 FILLER_27_24 ();
sky130_fd_sc_hd__decap_4 FILLER_27_3 ();
sky130_fd_sc_hd__decap_4 FILLER_27_31 ();
sky130_fd_sc_hd__decap_4 FILLER_27_38 ();
sky130_fd_sc_hd__decap_4 FILLER_27_45 ();
sky130_fd_sc_hd__decap_4 FILLER_27_52 ();
sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
sky130_fd_sc_hd__decap_8 FILLER_27_64 ();
sky130_fd_sc_hd__decap_12 FILLER_27_75 ();
sky130_fd_sc_hd__decap_4 FILLER_27_94 ();
sky130_fd_sc_hd__decap_6 FILLER_28_104 ();
sky130_fd_sc_hd__decap_8 FILLER_28_117 ();
sky130_fd_sc_hd__fill_2 FILLER_28_125 ();
sky130_fd_sc_hd__decap_6 FILLER_28_134 ();
sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
sky130_fd_sc_hd__decap_4 FILLER_28_15 ();
sky130_fd_sc_hd__decap_4 FILLER_28_150 ();
sky130_fd_sc_hd__decap_4 FILLER_28_161 ();
sky130_fd_sc_hd__decap_4 FILLER_28_168 ();
sky130_fd_sc_hd__decap_4 FILLER_28_175 ();
sky130_fd_sc_hd__fill_1 FILLER_28_179 ();
sky130_fd_sc_hd__decap_6 FILLER_28_187 ();
sky130_fd_sc_hd__fill_1 FILLER_28_19 ();
sky130_fd_sc_hd__fill_1 FILLER_28_193 ();
sky130_fd_sc_hd__decap_4 FILLER_28_23 ();
sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
sky130_fd_sc_hd__decap_3 FILLER_28_29 ();
sky130_fd_sc_hd__decap_6 FILLER_28_3 ();
sky130_fd_sc_hd__decap_4 FILLER_28_35 ();
sky130_fd_sc_hd__decap_4 FILLER_28_44 ();
sky130_fd_sc_hd__decap_12 FILLER_28_55 ();
sky130_fd_sc_hd__decap_4 FILLER_28_74 ();
sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
sky130_fd_sc_hd__decap_3 FILLER_28_85 ();
sky130_fd_sc_hd__decap_4 FILLER_28_93 ();
sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
sky130_fd_sc_hd__decap_12 FILLER_29_113 ();
sky130_fd_sc_hd__decap_4 FILLER_29_12 ();
sky130_fd_sc_hd__decap_8 FILLER_29_125 ();
sky130_fd_sc_hd__decap_3 FILLER_29_133 ();
sky130_fd_sc_hd__decap_8 FILLER_29_141 ();
sky130_fd_sc_hd__fill_1 FILLER_29_149 ();
sky130_fd_sc_hd__decap_6 FILLER_29_153 ();
sky130_fd_sc_hd__fill_1 FILLER_29_159 ();
sky130_fd_sc_hd__decap_4 FILLER_29_163 ();
sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
sky130_fd_sc_hd__decap_4 FILLER_29_178 ();
sky130_fd_sc_hd__decap_4 FILLER_29_189 ();
sky130_fd_sc_hd__fill_1 FILLER_29_193 ();
sky130_fd_sc_hd__decap_4 FILLER_29_21 ();
sky130_fd_sc_hd__fill_1 FILLER_29_25 ();
sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
sky130_fd_sc_hd__decap_4 FILLER_29_33 ();
sky130_fd_sc_hd__decap_6 FILLER_29_44 ();
sky130_fd_sc_hd__fill_1 FILLER_29_50 ();
sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
sky130_fd_sc_hd__decap_4 FILLER_29_66 ();
sky130_fd_sc_hd__fill_1 FILLER_29_70 ();
sky130_fd_sc_hd__decap_4 FILLER_29_78 ();
sky130_fd_sc_hd__decap_12 FILLER_29_87 ();
sky130_fd_sc_hd__decap_12 FILLER_29_99 ();
sky130_fd_sc_hd__decap_4 FILLER_2_110 ();
sky130_fd_sc_hd__decap_4 FILLER_2_117 ();
sky130_fd_sc_hd__fill_1 FILLER_2_121 ();
sky130_fd_sc_hd__decap_8 FILLER_2_129 ();
sky130_fd_sc_hd__decap_3 FILLER_2_137 ();
sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
sky130_fd_sc_hd__decap_6 FILLER_2_148 ();
sky130_fd_sc_hd__decap_12 FILLER_2_15 ();
sky130_fd_sc_hd__fill_1 FILLER_2_154 ();
sky130_fd_sc_hd__decap_4 FILLER_2_162 ();
sky130_fd_sc_hd__fill_1 FILLER_2_166 ();
sky130_fd_sc_hd__decap_8 FILLER_2_170 ();
sky130_fd_sc_hd__decap_4 FILLER_2_185 ();
sky130_fd_sc_hd__fill_2 FILLER_2_192 ();
sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
sky130_fd_sc_hd__decap_12 FILLER_2_29 ();
sky130_fd_sc_hd__decap_12 FILLER_2_3 ();
sky130_fd_sc_hd__fill_1 FILLER_2_41 ();
sky130_fd_sc_hd__decap_12 FILLER_2_49 ();
sky130_fd_sc_hd__decap_4 FILLER_2_61 ();
sky130_fd_sc_hd__decap_4 FILLER_2_72 ();
sky130_fd_sc_hd__fill_1 FILLER_2_76 ();
sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
sky130_fd_sc_hd__decap_6 FILLER_2_85 ();
sky130_fd_sc_hd__fill_1 FILLER_2_91 ();
sky130_fd_sc_hd__decap_4 FILLER_2_99 ();
sky130_fd_sc_hd__fill_1 FILLER_30_102 ();
sky130_fd_sc_hd__decap_12 FILLER_30_106 ();
sky130_fd_sc_hd__decap_4 FILLER_30_12 ();
sky130_fd_sc_hd__decap_12 FILLER_30_123 ();
sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
sky130_fd_sc_hd__decap_4 FILLER_30_146 ();
sky130_fd_sc_hd__decap_4 FILLER_30_155 ();
sky130_fd_sc_hd__decap_4 FILLER_30_166 ();
sky130_fd_sc_hd__decap_8 FILLER_30_173 ();
sky130_fd_sc_hd__fill_2 FILLER_30_181 ();
sky130_fd_sc_hd__decap_6 FILLER_30_188 ();
sky130_fd_sc_hd__decap_4 FILLER_30_23 ();
sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
sky130_fd_sc_hd__decap_6 FILLER_30_29 ();
sky130_fd_sc_hd__decap_6 FILLER_30_3 ();
sky130_fd_sc_hd__fill_1 FILLER_30_35 ();
sky130_fd_sc_hd__decap_4 FILLER_30_46 ();
sky130_fd_sc_hd__fill_1 FILLER_30_50 ();
sky130_fd_sc_hd__decap_4 FILLER_30_54 ();
sky130_fd_sc_hd__decap_4 FILLER_30_65 ();
sky130_fd_sc_hd__decap_12 FILLER_30_72 ();
sky130_fd_sc_hd__decap_4 FILLER_30_85 ();
sky130_fd_sc_hd__decap_6 FILLER_30_96 ();
sky130_fd_sc_hd__decap_6 FILLER_31_106 ();
sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
sky130_fd_sc_hd__decap_4 FILLER_31_122 ();
sky130_fd_sc_hd__decap_4 FILLER_31_13 ();
sky130_fd_sc_hd__decap_4 FILLER_31_133 ();
sky130_fd_sc_hd__decap_4 FILLER_31_144 ();
sky130_fd_sc_hd__decap_4 FILLER_31_155 ();
sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
sky130_fd_sc_hd__decap_4 FILLER_31_169 ();
sky130_fd_sc_hd__decap_4 FILLER_31_180 ();
sky130_fd_sc_hd__decap_3 FILLER_31_191 ();
sky130_fd_sc_hd__decap_4 FILLER_31_24 ();
sky130_fd_sc_hd__decap_3 FILLER_31_3 ();
sky130_fd_sc_hd__decap_4 FILLER_31_38 ();
sky130_fd_sc_hd__decap_4 FILLER_31_52 ();
sky130_fd_sc_hd__decap_4 FILLER_31_57 ();
sky130_fd_sc_hd__decap_4 FILLER_31_64 ();
sky130_fd_sc_hd__decap_4 FILLER_31_75 ();
sky130_fd_sc_hd__decap_4 FILLER_31_82 ();
sky130_fd_sc_hd__decap_6 FILLER_31_93 ();
sky130_fd_sc_hd__decap_6 FILLER_32_105 ();
sky130_fd_sc_hd__fill_1 FILLER_32_111 ();
sky130_fd_sc_hd__fill_2 FILLER_32_113 ();
sky130_fd_sc_hd__decap_4 FILLER_32_118 ();
sky130_fd_sc_hd__decap_4 FILLER_32_12 ();
sky130_fd_sc_hd__decap_4 FILLER_32_125 ();
sky130_fd_sc_hd__decap_8 FILLER_32_132 ();
sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
sky130_fd_sc_hd__decap_4 FILLER_32_146 ();
sky130_fd_sc_hd__decap_4 FILLER_32_153 ();
sky130_fd_sc_hd__decap_8 FILLER_32_160 ();
sky130_fd_sc_hd__fill_2 FILLER_32_169 ();
sky130_fd_sc_hd__decap_6 FILLER_32_174 ();
sky130_fd_sc_hd__decap_4 FILLER_32_190 ();
sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
sky130_fd_sc_hd__decap_4 FILLER_32_29 ();
sky130_fd_sc_hd__decap_6 FILLER_32_3 ();
sky130_fd_sc_hd__decap_4 FILLER_32_40 ();
sky130_fd_sc_hd__fill_2 FILLER_32_54 ();
sky130_fd_sc_hd__decap_8 FILLER_32_57 ();
sky130_fd_sc_hd__decap_4 FILLER_32_68 ();
sky130_fd_sc_hd__decap_4 FILLER_32_75 ();
sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
sky130_fd_sc_hd__decap_4 FILLER_32_90 ();
sky130_fd_sc_hd__fill_1 FILLER_32_94 ();
sky130_fd_sc_hd__decap_4 FILLER_32_98 ();
sky130_fd_sc_hd__decap_12 FILLER_3_100 ();
sky130_fd_sc_hd__decap_12 FILLER_3_113 ();
sky130_fd_sc_hd__decap_12 FILLER_3_125 ();
sky130_fd_sc_hd__decap_3 FILLER_3_137 ();
sky130_fd_sc_hd__decap_6 FILLER_3_143 ();
sky130_fd_sc_hd__decap_12 FILLER_3_15 ();
sky130_fd_sc_hd__decap_4 FILLER_3_152 ();
sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
sky130_fd_sc_hd__decap_4 FILLER_3_169 ();
sky130_fd_sc_hd__fill_1 FILLER_3_173 ();
sky130_fd_sc_hd__decap_4 FILLER_3_177 ();
sky130_fd_sc_hd__fill_1 FILLER_3_181 ();
sky130_fd_sc_hd__decap_4 FILLER_3_189 ();
sky130_fd_sc_hd__fill_1 FILLER_3_193 ();
sky130_fd_sc_hd__decap_8 FILLER_3_27 ();
sky130_fd_sc_hd__decap_12 FILLER_3_3 ();
sky130_fd_sc_hd__fill_1 FILLER_3_35 ();
sky130_fd_sc_hd__decap_4 FILLER_3_43 ();
sky130_fd_sc_hd__fill_1 FILLER_3_47 ();
sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
sky130_fd_sc_hd__decap_4 FILLER_3_57 ();
sky130_fd_sc_hd__fill_1 FILLER_3_61 ();
sky130_fd_sc_hd__decap_12 FILLER_3_65 ();
sky130_fd_sc_hd__decap_4 FILLER_3_77 ();
sky130_fd_sc_hd__fill_1 FILLER_3_81 ();
sky130_fd_sc_hd__decap_4 FILLER_3_85 ();
sky130_fd_sc_hd__fill_1 FILLER_3_89 ();
sky130_fd_sc_hd__decap_4 FILLER_3_93 ();
sky130_fd_sc_hd__decap_4 FILLER_4_101 ();
sky130_fd_sc_hd__fill_1 FILLER_4_105 ();
sky130_fd_sc_hd__decap_6 FILLER_4_111 ();
sky130_fd_sc_hd__fill_1 FILLER_4_117 ();
sky130_fd_sc_hd__decap_4 FILLER_4_125 ();
sky130_fd_sc_hd__decap_8 FILLER_4_132 ();
sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
sky130_fd_sc_hd__decap_4 FILLER_4_146 ();
sky130_fd_sc_hd__decap_12 FILLER_4_15 ();
sky130_fd_sc_hd__decap_4 FILLER_4_153 ();
sky130_fd_sc_hd__decap_8 FILLER_4_163 ();
sky130_fd_sc_hd__decap_4 FILLER_4_178 ();
sky130_fd_sc_hd__decap_4 FILLER_4_189 ();
sky130_fd_sc_hd__fill_1 FILLER_4_193 ();
sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
sky130_fd_sc_hd__decap_12 FILLER_4_3 ();
sky130_fd_sc_hd__decap_6 FILLER_4_35 ();
sky130_fd_sc_hd__decap_4 FILLER_4_48 ();
sky130_fd_sc_hd__decap_4 FILLER_4_55 ();
sky130_fd_sc_hd__fill_1 FILLER_4_59 ();
sky130_fd_sc_hd__decap_4 FILLER_4_66 ();
sky130_fd_sc_hd__decap_8 FILLER_4_73 ();
sky130_fd_sc_hd__decap_3 FILLER_4_81 ();
sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
sky130_fd_sc_hd__decap_6 FILLER_4_92 ();
sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
sky130_fd_sc_hd__decap_4 FILLER_5_113 ();
sky130_fd_sc_hd__decap_8 FILLER_5_124 ();
sky130_fd_sc_hd__fill_2 FILLER_5_132 ();
sky130_fd_sc_hd__decap_4 FILLER_5_141 ();
sky130_fd_sc_hd__decap_8 FILLER_5_150 ();
sky130_fd_sc_hd__decap_3 FILLER_5_165 ();
sky130_fd_sc_hd__decap_3 FILLER_5_169 ();
sky130_fd_sc_hd__fill_1 FILLER_5_17 ();
sky130_fd_sc_hd__fill_2 FILLER_5_192 ();
sky130_fd_sc_hd__decap_4 FILLER_5_25 ();
sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
sky130_fd_sc_hd__decap_8 FILLER_5_32 ();
sky130_fd_sc_hd__fill_1 FILLER_5_40 ();
sky130_fd_sc_hd__decap_4 FILLER_5_46 ();
sky130_fd_sc_hd__fill_1 FILLER_5_50 ();
sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
sky130_fd_sc_hd__decap_4 FILLER_5_66 ();
sky130_fd_sc_hd__decap_4 FILLER_5_77 ();
sky130_fd_sc_hd__decap_8 FILLER_5_88 ();
sky130_fd_sc_hd__decap_8 FILLER_5_9 ();
sky130_fd_sc_hd__fill_2 FILLER_5_96 ();
sky130_fd_sc_hd__fill_2 FILLER_6_100 ();
sky130_fd_sc_hd__decap_4 FILLER_6_105 ();
sky130_fd_sc_hd__fill_1 FILLER_6_109 ();
sky130_fd_sc_hd__decap_4 FILLER_6_116 ();
sky130_fd_sc_hd__decap_6 FILLER_6_12 ();
sky130_fd_sc_hd__decap_4 FILLER_6_123 ();
sky130_fd_sc_hd__decap_4 FILLER_6_130 ();
sky130_fd_sc_hd__decap_3 FILLER_6_137 ();
sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
sky130_fd_sc_hd__decap_6 FILLER_6_146 ();
sky130_fd_sc_hd__fill_1 FILLER_6_152 ();
sky130_fd_sc_hd__decap_6 FILLER_6_156 ();
sky130_fd_sc_hd__fill_1 FILLER_6_162 ();
sky130_fd_sc_hd__decap_4 FILLER_6_168 ();
sky130_fd_sc_hd__fill_1 FILLER_6_18 ();
sky130_fd_sc_hd__fill_2 FILLER_6_192 ();
sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
sky130_fd_sc_hd__decap_12 FILLER_6_36 ();
sky130_fd_sc_hd__decap_8 FILLER_6_51 ();
sky130_fd_sc_hd__fill_1 FILLER_6_59 ();
sky130_fd_sc_hd__decap_4 FILLER_6_63 ();
sky130_fd_sc_hd__decap_4 FILLER_6_70 ();
sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
sky130_fd_sc_hd__decap_4 FILLER_6_85 ();
sky130_fd_sc_hd__decap_8 FILLER_6_92 ();
sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
sky130_fd_sc_hd__decap_12 FILLER_7_113 ();
sky130_fd_sc_hd__decap_12 FILLER_7_125 ();
sky130_fd_sc_hd__decap_12 FILLER_7_137 ();
sky130_fd_sc_hd__decap_8 FILLER_7_149 ();
sky130_fd_sc_hd__fill_1 FILLER_7_15 ();
sky130_fd_sc_hd__fill_2 FILLER_7_157 ();
sky130_fd_sc_hd__decap_6 FILLER_7_162 ();
sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
sky130_fd_sc_hd__decap_3 FILLER_7_191 ();
sky130_fd_sc_hd__decap_12 FILLER_7_21 ();
sky130_fd_sc_hd__decap_12 FILLER_7_3 ();
sky130_fd_sc_hd__decap_3 FILLER_7_53 ();
sky130_fd_sc_hd__decap_8 FILLER_7_57 ();
sky130_fd_sc_hd__fill_1 FILLER_7_65 ();
sky130_fd_sc_hd__decap_4 FILLER_7_86 ();
sky130_fd_sc_hd__decap_12 FILLER_8_119 ();
sky130_fd_sc_hd__decap_4 FILLER_8_12 ();
sky130_fd_sc_hd__decap_8 FILLER_8_131 ();
sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
sky130_fd_sc_hd__decap_8 FILLER_8_163 ();
sky130_fd_sc_hd__fill_1 FILLER_8_171 ();
sky130_fd_sc_hd__fill_2 FILLER_8_192 ();
sky130_fd_sc_hd__decap_4 FILLER_8_23 ();
sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
sky130_fd_sc_hd__decap_4 FILLER_8_29 ();
sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
sky130_fd_sc_hd__fill_1 FILLER_8_33 ();
sky130_fd_sc_hd__decap_4 FILLER_8_54 ();
sky130_fd_sc_hd__decap_6 FILLER_8_78 ();
sky130_fd_sc_hd__decap_12 FILLER_8_85 ();
sky130_fd_sc_hd__fill_2 FILLER_8_97 ();
sky130_fd_sc_hd__decap_4 FILLER_9_107 ();
sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
sky130_fd_sc_hd__decap_4 FILLER_9_135 ();
sky130_fd_sc_hd__decap_8 FILLER_9_159 ();
sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
sky130_fd_sc_hd__decap_4 FILLER_9_18 ();
sky130_fd_sc_hd__decap_3 FILLER_9_191 ();
sky130_fd_sc_hd__decap_8 FILLER_9_25 ();
sky130_fd_sc_hd__decap_8 FILLER_9_3 ();
sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
sky130_fd_sc_hd__decap_8 FILLER_9_79 ();
sky130_fd_sc_hd__decap_3 PHY_0 ();
sky130_fd_sc_hd__decap_3 PHY_1 ();
sky130_fd_sc_hd__decap_3 PHY_10 ();
sky130_fd_sc_hd__decap_3 PHY_11 ();
sky130_fd_sc_hd__decap_3 PHY_12 ();
sky130_fd_sc_hd__decap_3 PHY_13 ();
sky130_fd_sc_hd__decap_3 PHY_14 ();
sky130_fd_sc_hd__decap_3 PHY_15 ();
sky130_fd_sc_hd__decap_3 PHY_16 ();
sky130_fd_sc_hd__decap_3 PHY_17 ();
sky130_fd_sc_hd__decap_3 PHY_18 ();
sky130_fd_sc_hd__decap_3 PHY_19 ();
sky130_fd_sc_hd__decap_3 PHY_2 ();
sky130_fd_sc_hd__decap_3 PHY_20 ();
sky130_fd_sc_hd__decap_3 PHY_21 ();
sky130_fd_sc_hd__decap_3 PHY_22 ();
sky130_fd_sc_hd__decap_3 PHY_23 ();
sky130_fd_sc_hd__decap_3 PHY_24 ();
sky130_fd_sc_hd__decap_3 PHY_25 ();
sky130_fd_sc_hd__decap_3 PHY_26 ();
sky130_fd_sc_hd__decap_3 PHY_27 ();
sky130_fd_sc_hd__decap_3 PHY_28 ();
sky130_fd_sc_hd__decap_3 PHY_29 ();
sky130_fd_sc_hd__decap_3 PHY_3 ();
sky130_fd_sc_hd__decap_3 PHY_30 ();
sky130_fd_sc_hd__decap_3 PHY_31 ();
sky130_fd_sc_hd__decap_3 PHY_32 ();
sky130_fd_sc_hd__decap_3 PHY_33 ();
sky130_fd_sc_hd__decap_3 PHY_34 ();
sky130_fd_sc_hd__decap_3 PHY_35 ();
sky130_fd_sc_hd__decap_3 PHY_36 ();
sky130_fd_sc_hd__decap_3 PHY_37 ();
sky130_fd_sc_hd__decap_3 PHY_38 ();
sky130_fd_sc_hd__decap_3 PHY_39 ();
sky130_fd_sc_hd__decap_3 PHY_4 ();
sky130_fd_sc_hd__decap_3 PHY_40 ();
sky130_fd_sc_hd__decap_3 PHY_41 ();
sky130_fd_sc_hd__decap_3 PHY_42 ();
sky130_fd_sc_hd__decap_3 PHY_43 ();
sky130_fd_sc_hd__decap_3 PHY_44 ();
sky130_fd_sc_hd__decap_3 PHY_45 ();
sky130_fd_sc_hd__decap_3 PHY_46 ();
sky130_fd_sc_hd__decap_3 PHY_47 ();
sky130_fd_sc_hd__decap_3 PHY_48 ();
sky130_fd_sc_hd__decap_3 PHY_49 ();
sky130_fd_sc_hd__decap_3 PHY_5 ();
sky130_fd_sc_hd__decap_3 PHY_50 ();
sky130_fd_sc_hd__decap_3 PHY_51 ();
sky130_fd_sc_hd__decap_3 PHY_52 ();
sky130_fd_sc_hd__decap_3 PHY_53 ();
sky130_fd_sc_hd__decap_3 PHY_54 ();
sky130_fd_sc_hd__decap_3 PHY_55 ();
sky130_fd_sc_hd__decap_3 PHY_56 ();
sky130_fd_sc_hd__decap_3 PHY_57 ();
sky130_fd_sc_hd__decap_3 PHY_58 ();
sky130_fd_sc_hd__decap_3 PHY_59 ();
sky130_fd_sc_hd__decap_3 PHY_6 ();
sky130_fd_sc_hd__decap_3 PHY_60 ();
sky130_fd_sc_hd__decap_3 PHY_61 ();
sky130_fd_sc_hd__decap_3 PHY_62 ();
sky130_fd_sc_hd__decap_3 PHY_63 ();
sky130_fd_sc_hd__decap_3 PHY_64 ();
sky130_fd_sc_hd__decap_3 PHY_65 ();
sky130_fd_sc_hd__decap_3 PHY_7 ();
sky130_fd_sc_hd__decap_3 PHY_8 ();
sky130_fd_sc_hd__decap_3 PHY_9 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
sky130_fd_sc_hd__clkbuf_4 _206_ (.A(net34),
.X(_097_));
sky130_fd_sc_hd__clkbuf_4 _207_ (.A(_097_),
.X(_098_));
sky130_fd_sc_hd__buf_2 _208_ (.A(_098_),
.X(_099_));
sky130_fd_sc_hd__xor2_1 _209_ (.A(\csa0.sc ),
.B(\csa0.y ),
.X(_100_));
sky130_fd_sc_hd__and2_1 _210_ (.A(\csa0.sc ),
.B(\csa0.y ),
.X(_101_));
sky130_fd_sc_hd__a31o_1 _211_ (.A1(_099_),
.A2(net2),
.A3(_100_),
.B1(_101_),
.X(_000_));
sky130_fd_sc_hd__nand2_1 _212_ (.A(_098_),
.B(net2),
.Y(_102_));
sky130_fd_sc_hd__xnor2_1 _213_ (.A(_102_),
.B(_100_),
.Y(\csa0.hsum2 ));
sky130_fd_sc_hd__a21o_1 _214_ (.A1(_097_),
.A2(net26),
.B1(\tcmp.z ),
.X(_032_));
sky130_fd_sc_hd__nand3_1 _215_ (.A(_097_),
.B(net26),
.C(\tcmp.z ),
.Y(_103_));
sky130_fd_sc_hd__and2_1 _216_ (.A(_032_),
.B(_103_),
.X(_104_));
sky130_fd_sc_hd__clkbuf_1 _217_ (.A(_104_),
.X(_031_));
sky130_fd_sc_hd__xor2_1 _218_ (.A(\genblk1[1].csa.sc ),
.B(\genblk1[1].csa.y ),
.X(_105_));
sky130_fd_sc_hd__and2_1 _219_ (.A(\genblk1[1].csa.sc ),
.B(\genblk1[1].csa.y ),
.X(_106_));
sky130_fd_sc_hd__a31o_1 _220_ (.A1(_099_),
.A2(net13),
.A3(_105_),
.B1(_106_),
.X(_011_));
sky130_fd_sc_hd__nand2_1 _221_ (.A(_098_),
.B(net13),
.Y(_107_));
sky130_fd_sc_hd__xnor2_1 _222_ (.A(_107_),
.B(_105_),
.Y(\genblk1[1].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _223_ (.A(\genblk1[2].csa.sc ),
.B(\genblk1[2].csa.y ),
.X(_108_));
sky130_fd_sc_hd__and2_1 _224_ (.A(\genblk1[2].csa.sc ),
.B(\genblk1[2].csa.y ),
.X(_109_));
sky130_fd_sc_hd__a31o_1 _225_ (.A1(_099_),
.A2(net24),
.A3(_108_),
.B1(_109_),
.X(_022_));
sky130_fd_sc_hd__nand2_1 _226_ (.A(_098_),
.B(net24),
.Y(_110_));
sky130_fd_sc_hd__xnor2_1 _227_ (.A(_110_),
.B(_108_),
.Y(\genblk1[2].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _228_ (.A(\genblk1[3].csa.sc ),
.B(\genblk1[3].csa.y ),
.X(_111_));
sky130_fd_sc_hd__and2_1 _229_ (.A(\genblk1[3].csa.sc ),
.B(\genblk1[3].csa.y ),
.X(_112_));
sky130_fd_sc_hd__a31o_1 _230_ (.A1(_099_),
.A2(net27),
.A3(_111_),
.B1(_112_),
.X(_024_));
sky130_fd_sc_hd__nand2_1 _231_ (.A(_098_),
.B(net27),
.Y(_113_));
sky130_fd_sc_hd__xnor2_1 _232_ (.A(_113_),
.B(_111_),
.Y(\genblk1[3].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _233_ (.A(\genblk1[4].csa.sc ),
.B(\genblk1[4].csa.y ),
.X(_114_));
sky130_fd_sc_hd__and2_1 _234_ (.A(\genblk1[4].csa.sc ),
.B(\genblk1[4].csa.y ),
.X(_115_));
sky130_fd_sc_hd__a31o_1 _235_ (.A1(_099_),
.A2(net28),
.A3(_114_),
.B1(_115_),
.X(_025_));
sky130_fd_sc_hd__nand2_1 _236_ (.A(_098_),
.B(net28),
.Y(_116_));
sky130_fd_sc_hd__xnor2_1 _237_ (.A(_116_),
.B(_114_),
.Y(\genblk1[4].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _238_ (.A(\genblk1[5].csa.sc ),
.B(\genblk1[5].csa.y ),
.X(_117_));
sky130_fd_sc_hd__and2_1 _239_ (.A(\genblk1[5].csa.sc ),
.B(\genblk1[5].csa.y ),
.X(_118_));
sky130_fd_sc_hd__a31o_1 _240_ (.A1(_099_),
.A2(net29),
.A3(_117_),
.B1(_118_),
.X(_026_));
sky130_fd_sc_hd__nand2_1 _241_ (.A(_098_),
.B(net29),
.Y(_119_));
sky130_fd_sc_hd__xnor2_1 _242_ (.A(_119_),
.B(_117_),
.Y(\genblk1[5].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _243_ (.A(\genblk1[6].csa.sc ),
.B(\genblk1[6].csa.y ),
.X(_120_));
sky130_fd_sc_hd__and2_1 _244_ (.A(\genblk1[6].csa.sc ),
.B(\genblk1[6].csa.y ),
.X(_121_));
sky130_fd_sc_hd__a31o_1 _245_ (.A1(_099_),
.A2(net30),
.A3(_120_),
.B1(_121_),
.X(_027_));
sky130_fd_sc_hd__clkbuf_4 _246_ (.A(_097_),
.X(_122_));
sky130_fd_sc_hd__nand2_1 _247_ (.A(_122_),
.B(net30),
.Y(_123_));
sky130_fd_sc_hd__xnor2_1 _248_ (.A(_123_),
.B(_120_),
.Y(\genblk1[6].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _249_ (.A(\genblk1[7].csa.sc ),
.B(\genblk1[7].csa.y ),
.X(_124_));
sky130_fd_sc_hd__and2_1 _250_ (.A(\genblk1[7].csa.sc ),
.B(\genblk1[7].csa.y ),
.X(_125_));
sky130_fd_sc_hd__a31o_1 _251_ (.A1(_099_),
.A2(net31),
.A3(_124_),
.B1(_125_),
.X(_028_));
sky130_fd_sc_hd__nand2_1 _252_ (.A(_122_),
.B(net31),
.Y(_126_));
sky130_fd_sc_hd__xnor2_1 _253_ (.A(_126_),
.B(_124_),
.Y(\genblk1[7].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _254_ (.A(\genblk1[8].csa.sc ),
.B(\genblk1[8].csa.y ),
.X(_127_));
sky130_fd_sc_hd__and2_1 _255_ (.A(\genblk1[8].csa.sc ),
.B(\genblk1[8].csa.y ),
.X(_128_));
sky130_fd_sc_hd__a31o_1 _256_ (.A1(_099_),
.A2(net32),
.A3(_127_),
.B1(_128_),
.X(_029_));
sky130_fd_sc_hd__nand2_1 _257_ (.A(_122_),
.B(net32),
.Y(_129_));
sky130_fd_sc_hd__xnor2_1 _258_ (.A(_129_),
.B(_127_),
.Y(\genblk1[8].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _259_ (.A(\genblk1[9].csa.sc ),
.B(\genblk1[10].csa.sum ),
.X(_130_));
sky130_fd_sc_hd__and2_1 _260_ (.A(\genblk1[9].csa.sc ),
.B(\genblk1[10].csa.sum ),
.X(_131_));
sky130_fd_sc_hd__a31o_1 _261_ (.A1(_099_),
.A2(net33),
.A3(_130_),
.B1(_131_),
.X(_030_));
sky130_fd_sc_hd__nand2_1 _262_ (.A(_122_),
.B(net33),
.Y(_132_));
sky130_fd_sc_hd__xnor2_1 _263_ (.A(_132_),
.B(_130_),
.Y(\genblk1[9].csa.hsum2 ));
sky130_fd_sc_hd__buf_2 _264_ (.A(_098_),
.X(_133_));
sky130_fd_sc_hd__xor2_1 _265_ (.A(\genblk1[10].csa.sc ),
.B(\genblk1[10].csa.y ),
.X(_134_));
sky130_fd_sc_hd__and2_1 _266_ (.A(\genblk1[10].csa.sc ),
.B(\genblk1[10].csa.y ),
.X(_135_));
sky130_fd_sc_hd__a31o_1 _267_ (.A1(_133_),
.A2(net3),
.A3(_134_),
.B1(_135_),
.X(_001_));
sky130_fd_sc_hd__nand2_1 _268_ (.A(_122_),
.B(net3),
.Y(_136_));
sky130_fd_sc_hd__xnor2_1 _269_ (.A(_136_),
.B(_134_),
.Y(\genblk1[10].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _270_ (.A(\genblk1[11].csa.sc ),
.B(\genblk1[11].csa.y ),
.X(_137_));
sky130_fd_sc_hd__and2_1 _271_ (.A(\genblk1[11].csa.sc ),
.B(\genblk1[11].csa.y ),
.X(_138_));
sky130_fd_sc_hd__a31o_1 _272_ (.A1(_133_),
.A2(net4),
.A3(_137_),
.B1(_138_),
.X(_002_));
sky130_fd_sc_hd__nand2_1 _273_ (.A(_122_),
.B(net4),
.Y(_139_));
sky130_fd_sc_hd__xnor2_1 _274_ (.A(_139_),
.B(_137_),
.Y(\genblk1[11].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _275_ (.A(\genblk1[12].csa.sc ),
.B(\genblk1[12].csa.y ),
.X(_140_));
sky130_fd_sc_hd__and2_1 _276_ (.A(\genblk1[12].csa.sc ),
.B(\genblk1[12].csa.y ),
.X(_141_));
sky130_fd_sc_hd__a31o_1 _277_ (.A1(_133_),
.A2(net5),
.A3(_140_),
.B1(_141_),
.X(_003_));
sky130_fd_sc_hd__nand2_1 _278_ (.A(_122_),
.B(net5),
.Y(_142_));
sky130_fd_sc_hd__xnor2_1 _279_ (.A(_142_),
.B(_140_),
.Y(\genblk1[12].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _280_ (.A(\genblk1[13].csa.sc ),
.B(\genblk1[13].csa.y ),
.X(_143_));
sky130_fd_sc_hd__and2_1 _281_ (.A(\genblk1[13].csa.sc ),
.B(\genblk1[13].csa.y ),
.X(_144_));
sky130_fd_sc_hd__a31o_1 _282_ (.A1(_133_),
.A2(net6),
.A3(_143_),
.B1(_144_),
.X(_004_));
sky130_fd_sc_hd__nand2_1 _283_ (.A(_122_),
.B(net6),
.Y(_145_));
sky130_fd_sc_hd__xnor2_1 _284_ (.A(_145_),
.B(_143_),
.Y(\genblk1[13].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _285_ (.A(\genblk1[14].csa.sc ),
.B(\genblk1[14].csa.y ),
.X(_146_));
sky130_fd_sc_hd__and2_1 _286_ (.A(\genblk1[14].csa.sc ),
.B(\genblk1[14].csa.y ),
.X(_147_));
sky130_fd_sc_hd__a31o_1 _287_ (.A1(_133_),
.A2(net7),
.A3(_146_),
.B1(_147_),
.X(_005_));
sky130_fd_sc_hd__nand2_1 _288_ (.A(_122_),
.B(net7),
.Y(_148_));
sky130_fd_sc_hd__xnor2_1 _289_ (.A(_148_),
.B(_146_),
.Y(\genblk1[14].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _290_ (.A(\genblk1[15].csa.sc ),
.B(\genblk1[15].csa.y ),
.X(_149_));
sky130_fd_sc_hd__and2_1 _291_ (.A(\genblk1[15].csa.sc ),
.B(\genblk1[15].csa.y ),
.X(_150_));
sky130_fd_sc_hd__a31o_1 _292_ (.A1(_133_),
.A2(net8),
.A3(_149_),
.B1(_150_),
.X(_006_));
sky130_fd_sc_hd__nand2_1 _293_ (.A(_122_),
.B(net8),
.Y(_151_));
sky130_fd_sc_hd__xnor2_1 _294_ (.A(_151_),
.B(_149_),
.Y(\genblk1[15].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _295_ (.A(\genblk1[16].csa.sc ),
.B(\genblk1[16].csa.y ),
.X(_152_));
sky130_fd_sc_hd__and2_1 _296_ (.A(\genblk1[16].csa.sc ),
.B(\genblk1[16].csa.y ),
.X(_153_));
sky130_fd_sc_hd__a31o_1 _297_ (.A1(_133_),
.A2(net9),
.A3(_152_),
.B1(_153_),
.X(_007_));
sky130_fd_sc_hd__buf_2 _298_ (.A(_097_),
.X(_154_));
sky130_fd_sc_hd__nand2_1 _299_ (.A(_154_),
.B(net9),
.Y(_155_));
sky130_fd_sc_hd__xnor2_1 _300_ (.A(_155_),
.B(_152_),
.Y(\genblk1[16].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _301_ (.A(\genblk1[17].csa.sc ),
.B(\genblk1[17].csa.y ),
.X(_156_));
sky130_fd_sc_hd__and2_1 _302_ (.A(\genblk1[17].csa.sc ),
.B(\genblk1[17].csa.y ),
.X(_157_));
sky130_fd_sc_hd__a31o_1 _303_ (.A1(_133_),
.A2(net10),
.A3(_156_),
.B1(_157_),
.X(_008_));
sky130_fd_sc_hd__nand2_1 _304_ (.A(_154_),
.B(net10),
.Y(_158_));
sky130_fd_sc_hd__xnor2_1 _305_ (.A(_158_),
.B(_156_),
.Y(\genblk1[17].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _306_ (.A(\genblk1[18].csa.sc ),
.B(\genblk1[18].csa.y ),
.X(_159_));
sky130_fd_sc_hd__and2_1 _307_ (.A(\genblk1[18].csa.sc ),
.B(\genblk1[18].csa.y ),
.X(_160_));
sky130_fd_sc_hd__a31o_1 _308_ (.A1(_133_),
.A2(net11),
.A3(_159_),
.B1(_160_),
.X(_009_));
sky130_fd_sc_hd__nand2_1 _309_ (.A(_154_),
.B(net11),
.Y(_161_));
sky130_fd_sc_hd__xnor2_1 _310_ (.A(_161_),
.B(_159_),
.Y(\genblk1[18].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _311_ (.A(\genblk1[19].csa.sc ),
.B(\genblk1[19].csa.y ),
.X(_162_));
sky130_fd_sc_hd__and2_1 _312_ (.A(\genblk1[19].csa.sc ),
.B(\genblk1[19].csa.y ),
.X(_163_));
sky130_fd_sc_hd__a31o_1 _313_ (.A1(_133_),
.A2(net12),
.A3(_162_),
.B1(_163_),
.X(_010_));
sky130_fd_sc_hd__nand2_1 _314_ (.A(_154_),
.B(net12),
.Y(_164_));
sky130_fd_sc_hd__xnor2_1 _315_ (.A(_164_),
.B(_162_),
.Y(\genblk1[19].csa.hsum2 ));
sky130_fd_sc_hd__clkbuf_4 _316_ (.A(_098_),
.X(_165_));
sky130_fd_sc_hd__xor2_1 _317_ (.A(\genblk1[20].csa.sc ),
.B(\genblk1[20].csa.y ),
.X(_166_));
sky130_fd_sc_hd__and2_1 _318_ (.A(\genblk1[20].csa.sc ),
.B(\genblk1[20].csa.y ),
.X(_167_));
sky130_fd_sc_hd__a31o_1 _319_ (.A1(_165_),
.A2(net14),
.A3(_166_),
.B1(_167_),
.X(_012_));
sky130_fd_sc_hd__nand2_1 _320_ (.A(_154_),
.B(net14),
.Y(_168_));
sky130_fd_sc_hd__xnor2_1 _321_ (.A(_168_),
.B(_166_),
.Y(\genblk1[20].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _322_ (.A(\genblk1[21].csa.sc ),
.B(\genblk1[21].csa.y ),
.X(_169_));
sky130_fd_sc_hd__and2_1 _323_ (.A(\genblk1[21].csa.sc ),
.B(\genblk1[21].csa.y ),
.X(_170_));
sky130_fd_sc_hd__a31o_1 _324_ (.A1(_165_),
.A2(net15),
.A3(_169_),
.B1(_170_),
.X(_013_));
sky130_fd_sc_hd__nand2_1 _325_ (.A(_154_),
.B(net15),
.Y(_171_));
sky130_fd_sc_hd__xnor2_1 _326_ (.A(_171_),
.B(_169_),
.Y(\genblk1[21].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _327_ (.A(\genblk1[22].csa.sc ),
.B(\genblk1[22].csa.y ),
.X(_172_));
sky130_fd_sc_hd__and2_1 _328_ (.A(\genblk1[22].csa.sc ),
.B(\genblk1[22].csa.y ),
.X(_173_));
sky130_fd_sc_hd__a31o_1 _329_ (.A1(_165_),
.A2(net16),
.A3(_172_),
.B1(_173_),
.X(_014_));
sky130_fd_sc_hd__nand2_1 _330_ (.A(_154_),
.B(net16),
.Y(_174_));
sky130_fd_sc_hd__xnor2_1 _331_ (.A(_174_),
.B(_172_),
.Y(\genblk1[22].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _332_ (.A(\genblk1[23].csa.sc ),
.B(\genblk1[23].csa.y ),
.X(_175_));
sky130_fd_sc_hd__and2_1 _333_ (.A(\genblk1[23].csa.sc ),
.B(\genblk1[23].csa.y ),
.X(_176_));
sky130_fd_sc_hd__a31o_1 _334_ (.A1(_165_),
.A2(net17),
.A3(_175_),
.B1(_176_),
.X(_015_));
sky130_fd_sc_hd__nand2_1 _335_ (.A(_154_),
.B(net17),
.Y(_177_));
sky130_fd_sc_hd__xnor2_1 _336_ (.A(_177_),
.B(_175_),
.Y(\genblk1[23].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _337_ (.A(\genblk1[24].csa.sc ),
.B(\genblk1[24].csa.y ),
.X(_178_));
sky130_fd_sc_hd__and2_1 _338_ (.A(\genblk1[24].csa.sc ),
.B(\genblk1[24].csa.y ),
.X(_179_));
sky130_fd_sc_hd__a31o_1 _339_ (.A1(_165_),
.A2(net18),
.A3(_178_),
.B1(_179_),
.X(_016_));
sky130_fd_sc_hd__nand2_1 _340_ (.A(_154_),
.B(net18),
.Y(_180_));
sky130_fd_sc_hd__xnor2_1 _341_ (.A(_180_),
.B(_178_),
.Y(\genblk1[24].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _342_ (.A(\genblk1[25].csa.sc ),
.B(\genblk1[25].csa.y ),
.X(_181_));
sky130_fd_sc_hd__and2_1 _343_ (.A(\genblk1[25].csa.sc ),
.B(\genblk1[25].csa.y ),
.X(_182_));
sky130_fd_sc_hd__a31o_1 _344_ (.A1(_165_),
.A2(net19),
.A3(_181_),
.B1(_182_),
.X(_017_));
sky130_fd_sc_hd__nand2_1 _345_ (.A(_154_),
.B(net19),
.Y(_183_));
sky130_fd_sc_hd__xnor2_1 _346_ (.A(_183_),
.B(_181_),
.Y(\genblk1[25].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _347_ (.A(\genblk1[26].csa.sc ),
.B(\genblk1[26].csa.y ),
.X(_184_));
sky130_fd_sc_hd__and2_1 _348_ (.A(\genblk1[26].csa.sc ),
.B(\genblk1[26].csa.y ),
.X(_185_));
sky130_fd_sc_hd__a31o_1 _349_ (.A1(_165_),
.A2(net20),
.A3(_184_),
.B1(_185_),
.X(_018_));
sky130_fd_sc_hd__nand2_1 _350_ (.A(_097_),
.B(net20),
.Y(_186_));
sky130_fd_sc_hd__xnor2_1 _351_ (.A(_186_),
.B(_184_),
.Y(\genblk1[26].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _352_ (.A(\genblk1[27].csa.sc ),
.B(\genblk1[27].csa.y ),
.X(_187_));
sky130_fd_sc_hd__and2_1 _353_ (.A(\genblk1[27].csa.sc ),
.B(\genblk1[27].csa.y ),
.X(_188_));
sky130_fd_sc_hd__a31o_1 _354_ (.A1(_165_),
.A2(net21),
.A3(_187_),
.B1(_188_),
.X(_019_));
sky130_fd_sc_hd__nand2_1 _355_ (.A(_097_),
.B(net21),
.Y(_189_));
sky130_fd_sc_hd__xnor2_1 _356_ (.A(_189_),
.B(_187_),
.Y(\genblk1[27].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _357_ (.A(\genblk1[28].csa.sc ),
.B(\genblk1[28].csa.y ),
.X(_190_));
sky130_fd_sc_hd__and2_1 _358_ (.A(\genblk1[28].csa.sc ),
.B(\genblk1[28].csa.y ),
.X(_191_));
sky130_fd_sc_hd__a31o_1 _359_ (.A1(_165_),
.A2(net22),
.A3(_190_),
.B1(_191_),
.X(_020_));
sky130_fd_sc_hd__nand2_1 _360_ (.A(_097_),
.B(net22),
.Y(_192_));
sky130_fd_sc_hd__xnor2_1 _361_ (.A(_192_),
.B(_190_),
.Y(\genblk1[28].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _362_ (.A(\genblk1[29].csa.sc ),
.B(\genblk1[29].csa.y ),
.X(_193_));
sky130_fd_sc_hd__and2_1 _363_ (.A(\genblk1[29].csa.sc ),
.B(\genblk1[29].csa.y ),
.X(_194_));
sky130_fd_sc_hd__a31o_1 _364_ (.A1(_165_),
.A2(net23),
.A3(_193_),
.B1(_194_),
.X(_021_));
sky130_fd_sc_hd__nand2_1 _365_ (.A(_097_),
.B(net23),
.Y(_195_));
sky130_fd_sc_hd__xnor2_1 _366_ (.A(_195_),
.B(_193_),
.Y(\genblk1[29].csa.hsum2 ));
sky130_fd_sc_hd__xor2_1 _367_ (.A(\genblk1[30].csa.sc ),
.B(\genblk1[30].csa.y ),
.X(_196_));
sky130_fd_sc_hd__and2_1 _368_ (.A(\genblk1[30].csa.sc ),
.B(\genblk1[30].csa.y ),
.X(_197_));
sky130_fd_sc_hd__a31o_1 _369_ (.A1(_098_),
.A2(net25),
.A3(_196_),
.B1(_197_),
.X(_023_));
sky130_fd_sc_hd__nand2_1 _370_ (.A(_097_),
.B(net25),
.Y(_198_));
sky130_fd_sc_hd__xnor2_1 _371_ (.A(_198_),
.B(_196_),
.Y(\genblk1[30].csa.hsum2 ));
sky130_fd_sc_hd__buf_4 _372_ (.A(net1),
.X(_199_));
sky130_fd_sc_hd__buf_4 _373_ (.A(_199_),
.X(_200_));
sky130_fd_sc_hd__inv_2 _374_ (.A(_200_),
.Y(_033_));
sky130_fd_sc_hd__inv_2 _375_ (.A(_200_),
.Y(_034_));
sky130_fd_sc_hd__inv_2 _376_ (.A(_200_),
.Y(_035_));
sky130_fd_sc_hd__inv_2 _377_ (.A(_200_),
.Y(_036_));
sky130_fd_sc_hd__inv_2 _378_ (.A(_200_),
.Y(_037_));
sky130_fd_sc_hd__inv_2 _379_ (.A(_200_),
.Y(_038_));
sky130_fd_sc_hd__inv_2 _380_ (.A(_200_),
.Y(_039_));
sky130_fd_sc_hd__inv_2 _381_ (.A(_200_),
.Y(_040_));
sky130_fd_sc_hd__inv_2 _382_ (.A(_200_),
.Y(_041_));
sky130_fd_sc_hd__inv_2 _383_ (.A(_200_),
.Y(_042_));
sky130_fd_sc_hd__buf_4 _384_ (.A(_199_),
.X(_201_));
sky130_fd_sc_hd__inv_2 _385_ (.A(_201_),
.Y(_043_));
sky130_fd_sc_hd__inv_2 _386_ (.A(_201_),
.Y(_044_));
sky130_fd_sc_hd__inv_2 _387_ (.A(_201_),
.Y(_045_));
sky130_fd_sc_hd__inv_2 _388_ (.A(_201_),
.Y(_046_));
sky130_fd_sc_hd__inv_2 _389_ (.A(_201_),
.Y(_047_));
sky130_fd_sc_hd__inv_2 _390_ (.A(_201_),
.Y(_048_));
sky130_fd_sc_hd__inv_2 _391_ (.A(_201_),
.Y(_049_));
sky130_fd_sc_hd__inv_2 _392_ (.A(_201_),
.Y(_050_));
sky130_fd_sc_hd__inv_2 _393_ (.A(_201_),
.Y(_051_));
sky130_fd_sc_hd__inv_2 _394_ (.A(_201_),
.Y(_052_));
sky130_fd_sc_hd__buf_4 _395_ (.A(_199_),
.X(_202_));
sky130_fd_sc_hd__inv_2 _396_ (.A(_202_),
.Y(_053_));
sky130_fd_sc_hd__inv_2 _397_ (.A(_202_),
.Y(_054_));
sky130_fd_sc_hd__inv_2 _398_ (.A(_202_),
.Y(_055_));
sky130_fd_sc_hd__inv_2 _399_ (.A(_202_),
.Y(_056_));
sky130_fd_sc_hd__inv_2 _400_ (.A(_202_),
.Y(_057_));
sky130_fd_sc_hd__inv_2 _401_ (.A(_202_),
.Y(_058_));
sky130_fd_sc_hd__inv_2 _402_ (.A(_202_),
.Y(_059_));
sky130_fd_sc_hd__inv_2 _403_ (.A(_202_),
.Y(_060_));
sky130_fd_sc_hd__inv_2 _404_ (.A(_202_),
.Y(_061_));
sky130_fd_sc_hd__inv_2 _405_ (.A(_202_),
.Y(_062_));
sky130_fd_sc_hd__buf_4 _406_ (.A(_199_),
.X(_203_));
sky130_fd_sc_hd__inv_2 _407_ (.A(_203_),
.Y(_063_));
sky130_fd_sc_hd__inv_2 _408_ (.A(_203_),
.Y(_064_));
sky130_fd_sc_hd__inv_2 _409_ (.A(_203_),
.Y(_065_));
sky130_fd_sc_hd__inv_2 _410_ (.A(_203_),
.Y(_066_));
sky130_fd_sc_hd__inv_2 _411_ (.A(_203_),
.Y(_067_));
sky130_fd_sc_hd__inv_2 _412_ (.A(_203_),
.Y(_068_));
sky130_fd_sc_hd__inv_2 _413_ (.A(_203_),
.Y(_069_));
sky130_fd_sc_hd__inv_2 _414_ (.A(_203_),
.Y(_070_));
sky130_fd_sc_hd__inv_2 _415_ (.A(_203_),
.Y(_071_));
sky130_fd_sc_hd__inv_2 _416_ (.A(_203_),
.Y(_072_));
sky130_fd_sc_hd__buf_4 _417_ (.A(_199_),
.X(_204_));
sky130_fd_sc_hd__inv_2 _418_ (.A(_204_),
.Y(_073_));
sky130_fd_sc_hd__inv_2 _419_ (.A(_204_),
.Y(_074_));
sky130_fd_sc_hd__inv_2 _420_ (.A(_204_),
.Y(_075_));
sky130_fd_sc_hd__inv_2 _421_ (.A(_204_),
.Y(_076_));
sky130_fd_sc_hd__inv_2 _422_ (.A(_204_),
.Y(_077_));
sky130_fd_sc_hd__inv_2 _423_ (.A(_204_),
.Y(_078_));
sky130_fd_sc_hd__inv_2 _424_ (.A(_204_),
.Y(_079_));
sky130_fd_sc_hd__inv_2 _425_ (.A(_204_),
.Y(_080_));
sky130_fd_sc_hd__inv_2 _426_ (.A(_204_),
.Y(_081_));
sky130_fd_sc_hd__inv_2 _427_ (.A(_204_),
.Y(_082_));
sky130_fd_sc_hd__buf_4 _428_ (.A(_199_),
.X(_205_));
sky130_fd_sc_hd__inv_2 _429_ (.A(_205_),
.Y(_083_));
sky130_fd_sc_hd__inv_2 _430_ (.A(_205_),
.Y(_084_));
sky130_fd_sc_hd__inv_2 _431_ (.A(_205_),
.Y(_085_));
sky130_fd_sc_hd__inv_2 _432_ (.A(_205_),
.Y(_086_));
sky130_fd_sc_hd__inv_2 _433_ (.A(_205_),
.Y(_087_));
sky130_fd_sc_hd__inv_2 _434_ (.A(_205_),
.Y(_088_));
sky130_fd_sc_hd__inv_2 _435_ (.A(_205_),
.Y(_089_));
sky130_fd_sc_hd__inv_2 _436_ (.A(_205_),
.Y(_090_));
sky130_fd_sc_hd__inv_2 _437_ (.A(_205_),
.Y(_091_));
sky130_fd_sc_hd__inv_2 _438_ (.A(_205_),
.Y(_092_));
sky130_fd_sc_hd__inv_2 _439_ (.A(_199_),
.Y(_093_));
sky130_fd_sc_hd__inv_2 _440_ (.A(_199_),
.Y(_094_));
sky130_fd_sc_hd__inv_2 _441_ (.A(_199_),
.Y(_095_));
sky130_fd_sc_hd__inv_2 _442_ (.A(_199_),
.Y(_096_));
sky130_fd_sc_hd__dfrtp_1 _443_ (.CLK(clknet_3_0__leaf_clk),
.D(_000_),
.RESET_B(_033_),
.Q(\csa0.sc ));
sky130_fd_sc_hd__dfrtp_1 _444_ (.CLK(clknet_3_1__leaf_clk),
.D(\csa0.hsum2 ),
.RESET_B(_034_),
.Q(net35));
sky130_fd_sc_hd__dfrtp_1 _445_ (.CLK(clknet_3_6__leaf_clk),
.D(_032_),
.RESET_B(_035_),
.Q(\tcmp.z ));
sky130_fd_sc_hd__dfrtp_1 _446_ (.CLK(clknet_3_4__leaf_clk),
.D(_031_),
.RESET_B(_036_),
.Q(\genblk1[30].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _447_ (.CLK(clknet_3_0__leaf_clk),
.D(_011_),
.RESET_B(_037_),
.Q(\genblk1[1].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _448_ (.CLK(clknet_3_1__leaf_clk),
.D(\genblk1[1].csa.hsum2 ),
.RESET_B(_038_),
.Q(\csa0.y ));
sky130_fd_sc_hd__dfrtp_1 _449_ (.CLK(clknet_3_0__leaf_clk),
.D(_022_),
.RESET_B(_039_),
.Q(\genblk1[2].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _450_ (.CLK(clknet_3_0__leaf_clk),
.D(\genblk1[2].csa.hsum2 ),
.RESET_B(_040_),
.Q(\genblk1[1].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _451_ (.CLK(clknet_3_1__leaf_clk),
.D(_024_),
.RESET_B(_041_),
.Q(\genblk1[3].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _452_ (.CLK(clknet_3_1__leaf_clk),
.D(\genblk1[3].csa.hsum2 ),
.RESET_B(_042_),
.Q(\genblk1[2].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _453_ (.CLK(clknet_3_0__leaf_clk),
.D(_025_),
.RESET_B(_043_),
.Q(\genblk1[4].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _454_ (.CLK(clknet_3_1__leaf_clk),
.D(\genblk1[4].csa.hsum2 ),
.RESET_B(_044_),
.Q(\genblk1[3].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _455_ (.CLK(clknet_3_1__leaf_clk),
.D(_026_),
.RESET_B(_045_),
.Q(\genblk1[5].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _456_ (.CLK(clknet_3_1__leaf_clk),
.D(\genblk1[5].csa.hsum2 ),
.RESET_B(_046_),
.Q(\genblk1[4].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _457_ (.CLK(clknet_3_4__leaf_clk),
.D(_027_),
.RESET_B(_047_),
.Q(\genblk1[6].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _458_ (.CLK(clknet_3_5__leaf_clk),
.D(\genblk1[6].csa.hsum2 ),
.RESET_B(_048_),
.Q(\genblk1[5].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _459_ (.CLK(clknet_3_4__leaf_clk),
.D(_028_),
.RESET_B(_049_),
.Q(\genblk1[7].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _460_ (.CLK(clknet_3_4__leaf_clk),
.D(\genblk1[7].csa.hsum2 ),
.RESET_B(_050_),
.Q(\genblk1[6].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _461_ (.CLK(clknet_3_0__leaf_clk),
.D(_029_),
.RESET_B(_051_),
.Q(\genblk1[8].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _462_ (.CLK(clknet_3_1__leaf_clk),
.D(\genblk1[8].csa.hsum2 ),
.RESET_B(_052_),
.Q(\genblk1[7].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _463_ (.CLK(clknet_3_0__leaf_clk),
.D(_030_),
.RESET_B(_053_),
.Q(\genblk1[9].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _464_ (.CLK(clknet_3_0__leaf_clk),
.D(\genblk1[9].csa.hsum2 ),
.RESET_B(_054_),
.Q(\genblk1[8].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _465_ (.CLK(clknet_3_2__leaf_clk),
.D(_001_),
.RESET_B(_055_),
.Q(\genblk1[10].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _466_ (.CLK(clknet_3_3__leaf_clk),
.D(\genblk1[10].csa.hsum2 ),
.RESET_B(_056_),
.Q(\genblk1[10].csa.sum ));
sky130_fd_sc_hd__dfrtp_1 _467_ (.CLK(clknet_3_2__leaf_clk),
.D(_002_),
.RESET_B(_057_),
.Q(\genblk1[11].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _468_ (.CLK(clknet_3_2__leaf_clk),
.D(\genblk1[11].csa.hsum2 ),
.RESET_B(_058_),
.Q(\genblk1[10].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _469_ (.CLK(clknet_3_2__leaf_clk),
.D(_003_),
.RESET_B(_059_),
.Q(\genblk1[12].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _470_ (.CLK(clknet_3_2__leaf_clk),
.D(\genblk1[12].csa.hsum2 ),
.RESET_B(_060_),
.Q(\genblk1[11].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _471_ (.CLK(clknet_3_2__leaf_clk),
.D(_004_),
.RESET_B(_061_),
.Q(\genblk1[13].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _472_ (.CLK(clknet_3_2__leaf_clk),
.D(\genblk1[13].csa.hsum2 ),
.RESET_B(_062_),
.Q(\genblk1[12].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _473_ (.CLK(clknet_3_2__leaf_clk),
.D(_005_),
.RESET_B(_063_),
.Q(\genblk1[14].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _474_ (.CLK(clknet_3_3__leaf_clk),
.D(\genblk1[14].csa.hsum2 ),
.RESET_B(_064_),
.Q(\genblk1[13].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _475_ (.CLK(clknet_3_6__leaf_clk),
.D(_006_),
.RESET_B(_065_),
.Q(\genblk1[15].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _476_ (.CLK(clknet_3_3__leaf_clk),
.D(\genblk1[15].csa.hsum2 ),
.RESET_B(_066_),
.Q(\genblk1[14].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _477_ (.CLK(clknet_3_3__leaf_clk),
.D(_007_),
.RESET_B(_067_),
.Q(\genblk1[16].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _478_ (.CLK(clknet_3_3__leaf_clk),
.D(\genblk1[16].csa.hsum2 ),
.RESET_B(_068_),
.Q(\genblk1[15].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _479_ (.CLK(clknet_3_2__leaf_clk),
.D(_008_),
.RESET_B(_069_),
.Q(\genblk1[17].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _480_ (.CLK(clknet_3_2__leaf_clk),
.D(\genblk1[17].csa.hsum2 ),
.RESET_B(_070_),
.Q(\genblk1[16].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _481_ (.CLK(clknet_3_3__leaf_clk),
.D(_009_),
.RESET_B(_071_),
.Q(\genblk1[18].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _482_ (.CLK(clknet_3_4__leaf_clk),
.D(\genblk1[18].csa.hsum2 ),
.RESET_B(_072_),
.Q(\genblk1[17].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _483_ (.CLK(clknet_3_3__leaf_clk),
.D(_010_),
.RESET_B(_073_),
.Q(\genblk1[19].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _484_ (.CLK(clknet_3_6__leaf_clk),
.D(\genblk1[19].csa.hsum2 ),
.RESET_B(_074_),
.Q(\genblk1[18].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _485_ (.CLK(clknet_3_6__leaf_clk),
.D(_012_),
.RESET_B(_075_),
.Q(\genblk1[20].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _486_ (.CLK(clknet_3_6__leaf_clk),
.D(\genblk1[20].csa.hsum2 ),
.RESET_B(_076_),
.Q(\genblk1[19].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _487_ (.CLK(clknet_3_6__leaf_clk),
.D(_013_),
.RESET_B(_077_),
.Q(\genblk1[21].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _488_ (.CLK(clknet_3_3__leaf_clk),
.D(\genblk1[21].csa.hsum2 ),
.RESET_B(_078_),
.Q(\genblk1[20].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _489_ (.CLK(clknet_3_6__leaf_clk),
.D(_014_),
.RESET_B(_079_),
.Q(\genblk1[22].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _490_ (.CLK(clknet_3_7__leaf_clk),
.D(\genblk1[22].csa.hsum2 ),
.RESET_B(_080_),
.Q(\genblk1[21].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _491_ (.CLK(clknet_3_7__leaf_clk),
.D(_015_),
.RESET_B(_081_),
.Q(\genblk1[23].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _492_ (.CLK(clknet_3_7__leaf_clk),
.D(\genblk1[23].csa.hsum2 ),
.RESET_B(_082_),
.Q(\genblk1[22].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _493_ (.CLK(clknet_3_5__leaf_clk),
.D(_016_),
.RESET_B(_083_),
.Q(\genblk1[24].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _494_ (.CLK(clknet_3_5__leaf_clk),
.D(\genblk1[24].csa.hsum2 ),
.RESET_B(_084_),
.Q(\genblk1[23].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _495_ (.CLK(clknet_3_7__leaf_clk),
.D(_017_),
.RESET_B(_085_),
.Q(\genblk1[25].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _496_ (.CLK(clknet_3_5__leaf_clk),
.D(\genblk1[25].csa.hsum2 ),
.RESET_B(_086_),
.Q(\genblk1[24].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _497_ (.CLK(clknet_3_7__leaf_clk),
.D(_018_),
.RESET_B(_087_),
.Q(\genblk1[26].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _498_ (.CLK(clknet_3_7__leaf_clk),
.D(\genblk1[26].csa.hsum2 ),
.RESET_B(_088_),
.Q(\genblk1[25].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _499_ (.CLK(clknet_3_7__leaf_clk),
.D(_019_),
.RESET_B(_089_),
.Q(\genblk1[27].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _500_ (.CLK(clknet_3_7__leaf_clk),
.D(\genblk1[27].csa.hsum2 ),
.RESET_B(_090_),
.Q(\genblk1[26].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _501_ (.CLK(clknet_3_5__leaf_clk),
.D(_020_),
.RESET_B(_091_),
.Q(\genblk1[28].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _502_ (.CLK(clknet_3_5__leaf_clk),
.D(\genblk1[28].csa.hsum2 ),
.RESET_B(_092_),
.Q(\genblk1[27].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _503_ (.CLK(clknet_3_5__leaf_clk),
.D(_021_),
.RESET_B(_093_),
.Q(\genblk1[29].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _504_ (.CLK(clknet_3_5__leaf_clk),
.D(\genblk1[29].csa.hsum2 ),
.RESET_B(_094_),
.Q(\genblk1[28].csa.y ));
sky130_fd_sc_hd__dfrtp_1 _505_ (.CLK(clknet_3_6__leaf_clk),
.D(_023_),
.RESET_B(_095_),
.Q(\genblk1[30].csa.sc ));
sky130_fd_sc_hd__dfrtp_1 _506_ (.CLK(clknet_3_4__leaf_clk),
.D(\genblk1[30].csa.hsum2 ),
.RESET_B(_096_),
.Q(\genblk1[29].csa.y ));
sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
.X(clknet_0_clk));
sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
.X(clknet_3_0__leaf_clk));
sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
.X(clknet_3_1__leaf_clk));
sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
.X(clknet_3_2__leaf_clk));
sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
.X(clknet_3_3__leaf_clk));
sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
.X(clknet_3_4__leaf_clk));
sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
.X(clknet_3_5__leaf_clk));
sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
.X(clknet_3_6__leaf_clk));
sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
.X(clknet_3_7__leaf_clk));
sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst),
.X(net1));
sky130_fd_sc_hd__clkbuf_1 input10 (.A(x[17]),
.X(net10));
sky130_fd_sc_hd__clkbuf_1 input11 (.A(x[18]),
.X(net11));
sky130_fd_sc_hd__clkbuf_1 input12 (.A(x[19]),
.X(net12));
sky130_fd_sc_hd__clkbuf_1 input13 (.A(x[1]),
.X(net13));
sky130_fd_sc_hd__clkbuf_1 input14 (.A(x[20]),
.X(net14));
sky130_fd_sc_hd__clkbuf_1 input15 (.A(x[21]),
.X(net15));
sky130_fd_sc_hd__clkbuf_1 input16 (.A(x[22]),
.X(net16));
sky130_fd_sc_hd__clkbuf_1 input17 (.A(x[23]),
.X(net17));
sky130_fd_sc_hd__clkbuf_1 input18 (.A(x[24]),
.X(net18));
sky130_fd_sc_hd__clkbuf_1 input19 (.A(x[25]),
.X(net19));
sky130_fd_sc_hd__clkbuf_1 input2 (.A(x[0]),
.X(net2));
sky130_fd_sc_hd__clkbuf_1 input20 (.A(x[26]),
.X(net20));
sky130_fd_sc_hd__clkbuf_1 input21 (.A(x[27]),
.X(net21));
sky130_fd_sc_hd__clkbuf_1 input22 (.A(x[28]),
.X(net22));
sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(x[29]),
.X(net23));
sky130_fd_sc_hd__clkbuf_1 input24 (.A(x[2]),
.X(net24));
sky130_fd_sc_hd__clkbuf_1 input25 (.A(x[30]),
.X(net25));
sky130_fd_sc_hd__clkbuf_1 input26 (.A(x[31]),
.X(net26));
sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(x[3]),
.X(net27));
sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(x[4]),
.X(net28));
sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(x[5]),
.X(net29));
sky130_fd_sc_hd__clkbuf_1 input3 (.A(x[10]),
.X(net3));
sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(x[6]),
.X(net30));
sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(x[7]),
.X(net31));
sky130_fd_sc_hd__clkbuf_1 input32 (.A(x[8]),
.X(net32));
sky130_fd_sc_hd__clkbuf_1 input33 (.A(x[9]),
.X(net33));
sky130_fd_sc_hd__clkbuf_1 input34 (.A(y),
.X(net34));
sky130_fd_sc_hd__clkbuf_1 input4 (.A(x[11]),
.X(net4));
sky130_fd_sc_hd__clkbuf_1 input5 (.A(x[12]),
.X(net5));
sky130_fd_sc_hd__clkbuf_1 input6 (.A(x[13]),
.X(net6));
sky130_fd_sc_hd__clkbuf_1 input7 (.A(x[14]),
.X(net7));
sky130_fd_sc_hd__clkbuf_1 input8 (.A(x[15]),
.X(net8));
sky130_fd_sc_hd__clkbuf_1 input9 (.A(x[16]),
.X(net9));
sky130_fd_sc_hd__buf_2 output35 (.A(net35),
.X(p));
endmodule
